module Exemplo(I1, I2, O)

input I1, I2;
output O;

and AND_1(O, I1, I2);

endmodule