module Exemplo(I1, I2, O1, O2);

input I1, I2;
output O1, O2;

and AND(O1, I1, I2);
or OR(O2, I1, I2);

endmodule